-- hello goiz this is our bery awn see-pee-you 
library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 